library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity hotelSystem_tb is
end entity hotelSystem_tb;

architecture rtl of hotelSystem_tb is
    
begin
    
    
    
end architecture rtl;